module mtc_ppa_mux_mpe #(
    parameter WIDTH_N = 2,//размер входного вектора request
    parameter AMOUNT_M = 1//максимальное число допустимых одновременных ответов
)(
    input   logic                                     clk,
    input   logic                                     reset_n,

    input   logic     [AMOUNT_M-1:0][WIDTH_N-1:0]     in_gnts_i,//th'
    input   logic     [AMOUNT_M-1:0][WIDTH_N-1:0]     in_gntss_i,//th''
    input   logic                                     in_gnt_vld_i,
    output  logic                                     in_gnt_rdy_o,

    output  logic     [AMOUNT_M-1:0][WIDTH_N-1:0]     out_gnt_o,
    output  logic                                     out_gnt_vld_o,
    input   logic                                     out_gnt_rdy_i
);

/***********************************************************************************************************************/
/***********************************************************************************************************************/
/*******************************************         DECLARATION         ***********************************************/
/***********************************************************************************************************************/
/***********************************************************************************************************************/
    logic [AMOUNT_M-1:0] selector;
    genvar i,j;

/***********************************************************************************************************************/
/***********************************************************************************************************************/
/*******************************************            LOGIC            ***********************************************/
/***********************************************************************************************************************/
/***********************************************************************************************************************/
    assign out_gnt_vld_o = in_gnt_vld_i;
    assign in_gnt_rdy_o = out_gnt_rdy_i;

    always_comb begin
        for(int i = 0; i < AMOUNT_M; i++) begin
            selector[i] = in_gnts_i[i][WIDTH_N-1];//нас интересуют только старшие биты
        end
    end


    generate
        //частный случай
        assign out_gnt_o[0] = selector[0] ? in_gnts_i[0] : in_gntss_i[0];

        for(i = 1; i < AMOUNT_M; i++) begin:gen_out_gnt//пробегаемся по всем массивам выходов
            //logic [0+:i][WIDTH_N-1:0] up_mux_out;//к глубокому сожалению динамический массив создать нельзя :-/
            logic [AMOUNT_M-1:0][WIDTH_N-1:0] up_mux_out;//к глубокому сожалению динамический массив создать нельзя :-/
            
            assign up_mux_out[0] = selector[0] ? in_gntss_i[i-1] : in_gntss_i[i];
            //а дальше пробегаемся по всем мультиплексорам
            for(j = 1; j <= i; j++)begin:gen_mux
                /*
                    i-j - для инвертирования порядка. Для того, чтобы понять как это работает - просто нарисуйте на бумаге и посмотрите :)
                */
                assign up_mux_out[j] = selector[j] ? ((j == i) ? in_gnts_i[j] : in_gntss_i[i-j-1]) : up_mux_out[j-1];//присваиваем значение из предыдущего мультиплексора в случае false
            end


            assign out_gnt_o[i] = up_mux_out[i];//присваиваем значение из последнего мультиплексора
        end
    endgenerate 

endmodule